*q3
V1 1 0 AC 1
R1 1 2 2k
R2 2 0 2k
C1 2 0 2u

.ac dec 100 1 20k
.end