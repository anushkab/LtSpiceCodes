*question 2
V1 1 0 PWL(0 12 0.001 24)
R1 1 2 4
L1 2 0 4
.tran 5
.end