*question 3
C1 1 0 0.1
R1 2 0 10
L1 1 2 1

.tran 4
.ic V(1,0)=10
.end