*question 1
C1 1 0 100u 
R2 1 2 1
R3 2 0 4
R4 2 0 4

.tran 1.5m
.ic V(1,0)=50
.end