*Question 3

V1 1 0 3
R1 1 2 10k
R2 2 0 15k
L1 2 0 3m

.tran 2

.end