* question 4
C1 1 0 4
R1 1 0 0.5
I1 0 1 10

.tran 10
.ic V(1,0)=2
.end