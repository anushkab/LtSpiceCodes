*q4
V1 1 0 AC sin(0 1 1)
C1 1 2 0.32u
Ra 2 3 10k
Rb 3 0 10k
C2 3 0 0.32u
R1 1 4 1k
R2 4 0 1k
.ac dec 100 1 100k
.end
