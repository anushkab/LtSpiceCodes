*q2
V1 1 0 AC sin(0 1 1)
C1 1 2 1u
R1 1 2 6k
R2 2 0 2k
.ac dec 100 1 1000
.end
 