*q3
V1 1 0 AC sin(0 1 1)
R1 1 2 40
L1 2 3 1.24m
C1 3 4 0.2u
C2 4 0 2u
R2 4 5 4
L2 5 0 0.124m
.ac dec 100 1 100k
.end