*q4
V1 1 0 AC 1
L1 1 2 0.0022
C1 2 3 47u
R1 3 0 13 
.ac dec 100 1 100k
.end