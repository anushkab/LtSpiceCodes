*question 2
V1 1 0 PWL(0 60 0.001 20)
R1 1 2 6
R2 2 0 3
C1 2 0 2

.tran 20
.end