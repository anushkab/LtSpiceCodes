*q1
I1 0 1 AC 1
C1 1 0 0.54p
R1 1 0 1k
L1 1 0 4u
.step param C1 0.54p 0.8p 0.1p
.ac dec 100 1 100M
.end