*question4

V1 1 0 PWL(0 10 1 10 1.001 0) 
R1 1 2 5
R2 2 0 20
L1 2 0 2

.tran 72
.end
